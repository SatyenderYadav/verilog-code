//////////////////////////////////////////////////////////////////////////////////
///////// [ SUM = A XOR B ] /////////////////////////////////////////////////////
///////// [ CARRY = A AND B ] //////////////////////////////////////////////////
module half_adder_data(a,b,sum,carry);
input a,b;
output sum,carry;

assign sum = a ^ b;
assign carry = a & b;
endmodule
/////////////////////////////////////////////////////////////////////////////////
///////// TEST BENCH ///////////////////////////////////////////////////////////
module half_adder_data_tb();
reg a,b;
wire sum,carry;
half_adder_data half_1(a,b,sum,carry);
initial
	begin
		a=0;b=0;
#10	a=0;b=1;
#10	a=1;b=0;
#10	a=1;b=1;
#10	
$stop;
end
endmodule
